* Equivalent circuit for state-space model from analysis of FastHenry file:
* * FastHenry2 File Automatically Generated.... JCCopyrights 2019

* Fasthenry generates  A dx/dt = x + B Vin,  Iout = C^t x + D Vin
* Note that regardless of what the original system modeled (say inductance),
* this file will use only R's, C's, and VCCS's to represent the system
* This is a 2-port model with the port nodes listed pairwise
* Correspondence to FastHenry nodes:
*   Port 1:  n66  to  n87, port name: secundary
*   Port 0:  n1  to  n65, port name: primary
* pn mn is a plus/minus port pair of nodes, where n is the port number

.subckt ROMequiv  p0 m0 p1 m1
* The coefficient of x is the identity == 1 ohm resistors to ground.
RH_0_0 state0 0 1
RH_1_1 state1 0 1
RH_2_2 state2 0 1
RH_3_3 state3 0 1

* The B matrix. VCCS dependent on port voltages
GB_0_0  state0 0 p0 m0         -1.2753
GB_1_1  state1 0 p1 m1        -2.12684
* The C matrix. VCCS dependent on state variable
GC_0_0   p0 m0 state0 0          1.2753
GC_1_1   p1 m1 state1 0         2.12684
GC_2_0   p0 m0 state2 0    1.40647e-013
GC_2_1   p1 m1 state2 0   -3.15737e-015
GC_3_0   p0 m0 state3 0    1.01715e-014
GC_3_1   p1 m1 state3 0     4.3319e-014
* The A matrix.  Coefficient of dx/dt.  constructed from capacitors. A = A^t
CA_0_0 state0 0   1.00345e-005 ic=0
CA_1_0 state1 state0  -2.58955e-007 ic=0
CA_1_1 state1 0   1.91961e-006 ic=0
CA_2_0 state2 state0   2.52667e-007 ic=0
CA_2_1 state2 state1    1.1199e-009 ic=0
CA_2_2 state2 0   8.73211e-008 ic=0
CA_3_1 state3 state1   4.90172e-008 ic=0
CA_3_2 state3 state2   2.25659e-010 ic=0
CA_3_3 state3 0   4.96677e-008 ic=0
.ends ROMequiv

* Equivalent circuit for state-space model from analysis of FastHenry file:
* * FastHenry2 File Automatically Generated.... JCCopyrights 2019

* Fasthenry generates  A dx/dt = x + B Vin,  Iout = C^t x + D Vin
* Note that regardless of what the original system modeled (say inductance),
* this file will use only R's, C's, and VCCS's to represent the system
* This is a 2-port model with the port nodes listed pairwise
* Correspondence to FastHenry nodes:
*   Port 1:  n126  to  n210, port name: secundary
*   Port 0:  n1  to  n125, port name: primary
* pn mn is a plus/minus port pair of nodes, where n is the port number

.subckt ROMequiv  p0 m0 p1 m1
* The coefficient of x is the identity == 1 ohm resistors to ground.
RH_0_0 state0 0 1
RH_1_1 state1 0 1
RH_2_2 state2 0 1
RH_3_3 state3 0 1

* The B matrix. VCCS dependent on port voltages
GB_0_0  state0 0 p0 m0        -7.94737
GB_1_1  state1 0 p1 m1        -5.64369
* The C matrix. VCCS dependent on state variable
GC_0_0   p0 m0 state0 0         7.94737
GC_1_1   p1 m1 state1 0         5.64369
GC_2_0   p0 m0 state2 0    6.28411e-013
GC_2_1   p1 m1 state2 0   -2.60804e-015
GC_3_0   p0 m0 state3 0     3.2205e-013
GC_3_1   p1 m1 state3 0    1.31946e-012
* The A matrix.  Coefficient of dx/dt.  constructed from capacitors. A = A^t
CA_0_0 state0 0    0.000394442 ic=0
CA_1_0 state1 state0  -5.30252e-006 ic=0
CA_1_1 state1 0   3.99323e-005 ic=0
CA_2_0 state2 state0   1.52329e-005 ic=0
CA_2_1 state2 state1   4.82438e-008 ic=0
CA_2_2 state2 0  -8.48612e-006 ic=0
CA_3_1 state3 state1   1.03438e-006 ic=0
CA_3_2 state3 state2   5.34186e-008 ic=0
CA_3_3 state3 0  -2.55635e-007 ic=0
.ends ROMequiv
